////////////////////////////////////////
// Company: Scaledge
// Engineer: Keertan Patel
// 
// Create Date: 4.5.2025 10:41:16
// Module Name: AHB_pkg
// Project Name: AHB slave verification 
// Description: pakage file
//
// v1.0 - File Created
///////////////////////////////////////


// guard statement to avoid multiple compilation of a file
`ifndef AHB_PKG_SV
`define AHB_PKG_SV

`include "AHB_defines.sv"
`include "AHB_inf.sv"

package AHB_pkg;
  `include "AHB_config.sv"
  `include "AHB_trans.sv"
  `include "AHB_gen.sv"
  `include "AHB_driver.sv"
  `include "AHB_mon.sv"
  `include "AHB_ref_model.sv"
  `include "AHB_scb.sv"
  `include "AHB_env.sv"
  `include "AHB_write_read.sv"
  `include "AHB_back_to_back.sv"
  `include "AHB_idle_test.sv"
  `include "AHB_base_test.sv"

 endpackage
`endif
