/*  -----------to do in driver file--------------
	
*/

/*-------------to do in generator file---------------
	-->create a queue named haddr_que and push all the addresses required for the transaction in it. it will be popped in driver.
*/